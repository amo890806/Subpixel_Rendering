`define HEADER 54
`define WIDTH 1080
`define HEIGHT 1920

`define HD 270      //HACT
`define HS 1       //HSYNC
`define HB 64       //HBP
`define HF 26       //HFP
`define HT 361      //HTOTAL
`define VD 1920     //HEIGHT / VACT
`define VS 1        //VSYNC
`define VB 33       //VBP
`define VF 10       //VFP
`define VT 1964     //VTOTAL

`define SHP_64 64*16
`define SHP_128 128*16
`define SHP_192 192*16
`define SHP_256 256*16
`define SPR_SHARP_amout 4*16

`define SPR_THR_B_edge 64
`define SPR_THR_R_edge 64

